* /home/win/working/cdi-tach/tach_pulse_sim/tach_pulse_filter.cir

* EESchema Netlist Version 1.1 (Spice format) creation date: Tue 11 Aug 2015 06:21:39 PM PDT

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

* Sheet Name: /
C1  0 TACH_OUT 22nF
R1  TACH_IN TACH_OUT 100K
R2  TACH_OUT 0 12.1K
*V1 TACH_IN 0 sin(0 40 50) dc=0 ac=10
V1 TACH_IN 0 pulse(0 40 0 1us 1us 4ms 8ms) dc=0 ac=1

.control
tran 1us 20ms
plot TACH_IN TACH_OUT
.endc
.end
